* /home/janakiram.emani/janakiram_elevator/elevator/elevator.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Fri 04 Mar 2022 08:00:12 AM UTC

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  ? ? ? ? ? ? ? ? ? janakiram_elevator		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U2-Pad7_ Net-_U2-Pad8_ Net-_U2-Pad9_ janakiram_elevator		
U3  clk0 rst0 ra0 rb0 rc0 rd0 Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ adc_bridge_6		
U4  Net-_U2-Pad7_ Net-_U2-Pad8_ Net-_U2-Pad9_ Net-_R1-Pad1_ Net-_R2-Pad1_ Net-_R3-Pad1_ dac_bridge_3		
v7  rd0 GND pulse		
v6  rc0 GND pulse		
v5  rb0 GND pulse		
v4  ra0 GND pulse		
v3  rst0 GND pulse		
v2  clk0 GND pulse		
R1  Net-_R1-Pad1_ floor1 1k		
R2  Net-_R2-Pad1_ floor0 1k		
R3  Net-_R3-Pad1_ dir0 1k		
C1  floor1 GND 1u		
C2  floor0 GND 1u		
C3  dir0 GND 1u		
U12  floor0 plot_v1		
U11  floor1 plot_v1		
U13  dir0 plot_v1		
U5  clk0 plot_v1		
U6  rst0 plot_v1		
U7  ra0 plot_v1		
U8  rb0 plot_v1		
U9  rc0 plot_v1		
U10  rd0 plot_v1		

.end
